function void fxn(int var1, var2);
  $display(var1, var2);
endfunction: fxn

function int product(input int var1, var2, output var3);
    product = var1 * var2;
    var3 = product*2;
endfunction
