module example();                                                   
    reg clock, reset, enable, data;                           

    initial                                                    
        begin
             clock = 0;                                     
             reset = 0;
             enable = 0;
             data = 0;
        end
endmodule
