module array();
  bit[7:0][7:0]bytes;
  $displayh(bytes,
    bytes[7],
    bytes[7][7]
  );
endmodule
