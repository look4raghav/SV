program test(temp_if intf);
  initial
    begin
      run();
    end
  task run ();
    a = RAGHAV
      $display("A = %d", a);
  endtask: run
endprogram: test
