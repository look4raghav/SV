module final_exp; 
    initial 
        #100 $finish; 
        final 
             $display(" END OF SIMULATION at %d ",$time); 
endmodule 
