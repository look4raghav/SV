class training_c;
  int coutse_fee;
  
function int total_subjects;
  return course_fee;
endfunction
endclass

Training_c train_h = new;
