Class training_c;
int coutse_fee;
function int total_subjects;
  return course_fee;
endfunction

task deposit(input int tax);
  course_fee = course_fee + tax;
endtask
endclass
