module array();
  int count, total, n[] = {1,4,6,15,8,3,10,05,16,12};
  
  count = n.sum with ((item > 7));
  total = n.sum with ((item < 7));
  
  n.reverse();
  n.sort();
  n.shuffle();
  n.rsort();
  
endmodule
